library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library work;
use work.cpu_defs.all;
use work.utils_pak.all;


entity controller_tb is end;

architecture controller_tb_arc of controller_tb is

    signal clk:             std_logic := '0';
    signal reset_n:         std_logic;
    signal mem_read:        std_logic;
    signal mem_write:       std_logic;
    signal mem_bytesel:     std_logic_vector(3 downto 0);
    signal mem_addr:        word;
    signal mem_data_out:    word;
    signal mem_ack:         std_logic;
    signal mem_data_in:     word;
    signal reg_sel_a:       std_logic_vector(4 downto 0);
    signal reg_a_out:       word;
    signal reg_sel_b:       std_logic_vector(4 downto 0);
    signal reg_b_out:       word;
    signal reg_sel_c:       std_logic_vector(4 downto 0);
    signal reg_c_out:       word;
    signal reg_sel_y:       std_logic_vector(4 downto 0);
    signal reg_write_y:     std_logic;
    signal reg_y_in:        word;
    signal reg_sel_z:       std_logic_vector(4 downto 0);
    signal reg_write_z:     std_logic;
    signal reg_z_in:        word;
    signal alu_op:          cpu_opcode;
    signal alu_rs_in:       word;
    signal alu_rt_in:       word;
    signal alu_rd_in:       word;
    signal alu_imm_in:      word;
    signal alu_output_a:    word;
    signal alu_output_b:    word;
    signal pc_in:           word;
    signal pc_write:        std_logic;
    signal pc_out:          word;
    signal dummy:           std_logic;

begin
    clk <= not clk after 14 ns;
    reset_n <= '0', '1' after 100 ns;

    -- Providing the controller with data from the memory.
    -- Simulating a synchronous memory read access
    --
    proc_mem_data_in: process(clk, reset_n)
    begin
        if (reset_n = '0') then
            mem_data_in <= (others => '0');
        elsif (rising_edge(clk)) then
            if mem_read = '1' then
                -- The reset address, provide first instruction
                if mem_addr = x"00100000" then
                    --
                    -- sub $r5, $r6, $r9
                    --
                    -- generated by luz_asm_sim test_assembler.py
                    --
                    mem_data_in <= x"04a64800";
                elsif mem_addr = x"00100004" then
                    --
                    -- mulu $r20, $r2, $r3
                    --
                    mem_data_in <= x"0A821800";
                end if;
            end if;
        end if;
    end process;
    
    -- Simulate the way the acknowledge signal from memory behaves
    --
    mem_ack <= '1' when mem_read = '1' or mem_write = '1' else '0';
    
    -- Simulate reading from register A (Rd)
    --
    proc_reg_a_out: process(clk, reset_n)
    begin
        if (reset_n = '0') then
            reg_a_out <= (others => '0');
        elsif (rising_edge(clk)) then
            if to_integer(unsigned(reg_sel_a)) = 6 then 
                reg_a_out <= x"0034AABB";
            else
                reg_a_out <= (others => '0');
            end if;
        end if;
    end process;

    -- Simulate reading from register B (Rs)
    --
    proc_reg_b_out: process(clk, reset_n)
    begin
        if (reset_n = '0') then
            reg_b_out <= (others => '0');
        elsif (rising_edge(clk)) then
            if to_integer(unsigned(reg_sel_b)) = 6 then 
                reg_b_out <= x"0034AABB";
            elsif to_integer(unsigned(reg_sel_b)) = 2 then 
                reg_b_out <= x"00400000";
            else
                reg_b_out <= (others => '0');
            end if;
        end if;
    end process;

    -- Simulate reading from register C (Rt)
    --
    proc_reg_c_out: process(clk, reset_n)
    begin
        if (reset_n = '0') then
            reg_c_out <= (others => '0');
        elsif (rising_edge(clk)) then
            if to_integer(unsigned(reg_sel_c)) = 9 then 
                reg_c_out <= x"00126789";
            elsif to_integer(unsigned(reg_sel_c)) = 3 then 
                reg_c_out <= x"00AB0000";
            else
                reg_c_out <= (others => '0');
            end if;
        end if;
    end process;


    process
    begin
        
        wait;
    end process;

    dut: entity work.controller(controller_arc)
    port map
    (
        clk             => clk,
        reset_n         => reset_n,
        mem_read        => mem_read,
        mem_write       => mem_write,
        mem_bytesel     => mem_bytesel,
        mem_addr        => mem_addr,
        mem_data_out    => mem_data_out,
        mem_ack         => mem_ack,
        mem_data_in     => mem_data_in,
        reg_sel_a       => reg_sel_a,
        reg_a_out       => reg_a_out,
        reg_sel_b       => reg_sel_b,
        reg_b_out       => reg_b_out,
        reg_sel_c       => reg_sel_c,
        reg_c_out       => reg_c_out,
        reg_sel_y       => reg_sel_y,
        reg_write_y     => reg_write_y,
        reg_y_in        => reg_y_in,
        reg_sel_z       => reg_sel_z,
        reg_write_z     => reg_write_z,
        reg_z_in        => reg_z_in,
        alu_op          => alu_op,
        alu_rs_in       => alu_rs_in,
        alu_rt_in       => alu_rt_in,
        alu_rd_in       => alu_rd_in,
        alu_imm_in      => alu_imm_in,
        alu_output_a    => alu_output_a,
        alu_output_b    => alu_output_b,
        pc_in           => pc_in,
        pc_write        => pc_write,
        pc_out          => pc_out,
        dummy           => dummy
    );
    
    pc_map: entity work.program_counter(program_counter_arc)
    generic map
    (
        INIT        => x"00100000"
    )
    port map
    (
        clk         => clk,
        reset_n     => reset_n,
        pc_in       => pc_in,
        pc_out      => pc_out,
        pc_write    => pc_write
    );
    
    alu_map: entity work.alu(alu_arc)
    port map
    (
        clk         => clk,
        reset_n     => reset_n,
        op          => alu_op,
        rd_in       => alu_rd_in,
        rt_in       => alu_rt_in,
        rs_in       => alu_rs_in,
        imm_in      => alu_imm_in,
        output_a    => alu_output_a,
        output_b    => alu_output_b
    );
    
end;

